/*
 * Copyright (c) 2025 Matthew Chen, Jovan Koledin, Ryan Leahy
 * SPDX-License-Identifier: Apache-2.0
 */

module vga (
    output reg [9:0] vaddr,
    output reg [9:0] haddr,
    output reg vsync,
    output reg hsync,

    input wire rst,
    input wire clk
);


endmodule